----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    20:39:52 09/12/2018 
-- Design Name: 
-- Module Name:    nibble7seg - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity nibble7seg is
    Port ( selectionEntry : in  STD_LOGIC_VECTOR (7 downto 0);
           nibbleOutputLSN : out  STD_LOGIC_VECTOR (6 downto 0);
			  nibbleOutputMSN : out  STD_LOGIC_VECTOR (6 downto 0));
end nibble7seg;

architecture Behavioral of nibble7seg is
	signal msN : STD_LOGIC_VECTOR (6 downto 0);
	signal lsN : STD_LOGIC_VECTOR (6 downto 0);
begin
	with selectionEntry(7 downto 4) select
		msN <= 	"0000001" when "0000", -- '0'
					"1001111" when "0001", -- '1'
					"0010010" when "0010", -- '2'
					"0000110" when "0011", -- '3'
					"1001100" when "0100", -- '4'
					"0100100" when "0101", -- '5'
					"0100000" when "0110", -- '6'
					"0001111" when "0111", -- '7'
					"0000000" when "1000", -- '8'
					"0000100" when "1001", -- '9'
					"0001000" when "1010", -- 'A'
					"1100000" when "1011", -- 'B'
					"0110001" when "1100", -- 'C'
					"1000010" when "1101", -- 'D'
					"0110000" when "1110", -- 'E'
					"0111000" when "1111", -- 'F'
					"1111111" when others;
	
	with selectionEntry(3 downto 0) select
		lsN <=	"0000001" when "0000", -- '0'
					"1001111" when "0001", -- '1'
					"0010010" when "0010", -- '2'
					"0000110" when "0011", -- '3'
					"1001100" when "0100", -- '4'
					"0100100" when "0101", -- '5'
					"0100000" when "0110", -- '6'
					"0001111" when "0111", -- '7'
					"0000000" when "1000", -- '8'
					"0000100" when "1001", -- '9'
					"0001000" when "1010", -- 'A'
					"1100000" when "1011", -- 'B'
					"0110001" when "1100", -- 'C'
					"1000010" when "1101", -- 'D'
					"0110000" when "1110", -- 'E'
					"0111000" when "1111", -- 'F'
					"1111111" when others;

	nibbleOutputMSN(6 downto 0) <= msN;
	nibbleOutputLSN(6 downto 0) <= lsN;
end Behavioral;

